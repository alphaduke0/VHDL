force sim:/mux4x1/E 1010;
run;

force sim:/mux4x1/S 01; run;
force sim:/mux4x1/S 10; run;
force sim:/mux4x1/S 11; run;
force sim:/mux4x1/S 00; run;